netcdf sres-a1b_ukcp18-land-prob-25km_sample_day_19981201-19991130 {
dimensions:
	time = 2 ;
	lat = 2 ;
	lon = 2 ;
variables:
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "Time" ;
		time:axis = "T" ;
		time:units = "seconds since 1970-01-01T00:00:00Z" ;
	float lat ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:axis = "Y" ;
		lat:long_name = "Latitude" ;
	float lon ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:axis = "X" ;
		lon:long_name = "Longitude" ;
	float z ;
		z:standard_name = "depth" ;
		z:positive = "down" ;
		z:units = "m" ;
		z:long_name = "Depth below surface" ;
	float temperature(time, lat, lon) ;
		temperature:standard_name = "sea_water_temperature" ;
		temperature:units = "deg_C" ;
		temperature:long_name = "Seawater Temperature" ;
		temperature:coordinates = "time lat lon z" ;

// global attributes:
		:Conventions = "CF-1.5" ;
		:variable = "tas" ;
		:scenario = "sres-a1b" ;
		:prob_data_type = "sample" ;
		:dataset_id = "ukcp18-land-prob-25km" ;
		:frequency = "day" ;
data:

 time = _, _ ;

 lat = _ ;

 lon = _ ;

 z = _ ;

 temperature =
  _, _,
  _, _,
  _, _,
  _, _ ;
}

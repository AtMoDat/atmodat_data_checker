netcdf simple_nc4 {
dimensions:
	time = 2 ;
	lat = 2 ;
	lon = 2 ;
variables:
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "Time" ;
		time:axis = "T" ;
		time:units = "seconds since 1970-01-01T00:00:00Z" ;
	float lat(lat);
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:axis = "Y" ;
		lat:long_name = "Latitude" ;
	float lon(lon);
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:axis = "X" ;
		lon:long_name = "Longitude" ;
	float z ;
		z:standard_name = "depth" ;
		z:positive = "down" ;
		z:units = "m" ;
		z:long_name = "Depth below surface" ;
	float temperature(time, lat, lon) ;
		temperature:standard_name = "sea_water_temperature" ;
		temperature:units = "deg_C" ;
		temperature:long_name = "Seawater Temperature" ;
		temperature:coordinates = "time lat lon z" ;

// global attributes:
		:Conventions = "CF-1.5" ;
		:source = "Good data from a good place." ;
		:project_id = "EUSTACE" ;
		:contact = "My name, my address." ;
		:history = "Created in the past by people." ;
		:references = "Wilson, A.B.C. (1999). Etc" ;
		:product_version = "MERIS X.Y" ;
		:title = "A very splendid data product" ;
		:summary = "A very very very splendid data product." ;
		:creator_name = "Mrs Brilliant" ;
		:creator_email = "mrs.brilliant@the.world" ;
		:frequency = "day" ;
		:institution_id = "MOHC" ;
		:institution = "Met Office Hadley Centre, Fitzroy Road, Exeter, Devon, EX1 3PB, UK" ;
		:creation_date = "2020-01-20T20:20:20" ;
data:

 time = 100, 101 ;

 lat = 20 ;

 lon = 40 ;

 z = 1 ;

 temperature =
  21, 23,
  12, 34,
  8, 16,
  18, 19 ;
}

netcdf tasAnom_rcp85_land-prob_uk_25km_cdf_mon_20001201-20011130 {
dimensions:
	percentile = 111 ;
	projection_x_coordinate = 1 ;
	projection_y_coordinate = 2 ;
	time = UNLIMITED ; // (0 currently)
variables:
	double percentile(percentile) ;
		percentile:long_name = "percentile" ;
	double projection_x_coordinate(projection_x_coordinate) ;
		projection_x_coordinate:units = "m" ;
		projection_x_coordinate:standard_name = "projection_x_coordinate" ;
		projection_x_coordinate:bounds = "projection_x_coordinate_bnds" ;
		projection_x_coordinate:axis = "X" ;
	double projection_y_coordinate(projection_y_coordinate) ;
		projection_y_coordinate:units = "m" ;
		projection_y_coordinate:standard_name = "projection_y_coordinate" ;
		projection_y_coordinate:bounds = "projection_y_coordinate_bnds" ;
		projection_y_coordinate:axis = "Y" ;
	float tasAnom(time, projection_y_coordinate, projection_x_coordinate, percentile) ;
		tasAnom:_FillValue = 1.e+20f ;
		tasAnom:anomaly_type = "absolute_change" ;
		tasAnom:grid_mapping = "transverse_mercator" ;
		tasAnom:description = "Surface temperature anomaly at 1.5m (°c)" ;
		tasAnom:baseline_period = "1981-2000" ;
		tasAnom:coordinates = "latitude longitude season_year" ;
		tasAnom:long_name = "Anomaly of air temperature" ;
		tasAnom:standard_name = "air_temperature" ;
		tasAnom:cell_methods = "time: mean" ;
		tasAnom:units = "K" ;
	float time(time) ;
		time:units = "days since 2000-12-15 00:00:00" ;
		time:long_name = "Time" ;
		time:calendar = "360_day" ;
		time:standard_name = "time" ;
		time:bounds = "time_bounds" ;

// global attributes:
		:variable = "tasAnom" ;
		:institution_id = "MOHC" ;
		:domain = "uk" ;
		:scenario = "rcp85" ;
		:creator_name = "***Your name***" ;
		:title = "***Title of my data set***" ;
		:creator_email = "***Your email***" ;
		:baseline_period = "1981-2000" ;
		:institution = "Met Office Hadley Centre (MOHC), FitzRoy Road, Exeter, Devon, EX1 3PB, UK." ;
		:collection = "land-prob" ;
		:creation_date = "2018-03-31 12:00:00" ;
		:project = "ukcp18" ;
		:source = "***The method of production of the original data. If it was model-generated, source should name the model and its version, as specifically as could be useful.***" ;
		:frequency = "mon" ;
		:references = "https://www.metoffice.gov.uk/***NEW**UKCP**SITE***" ;
		:contact = "***Required from Fai***" ;
		:version = "v20180331" ;
		:dataset_id = "ukcp18-land-prob-uk-25km-all" ;
		:resolution = "25km" ;
		:prob_data_type = "cdf" ;
		:history = "Tue Mar 20 14:35:49 2018: ncks -d projection_y_coordinate,,,50 -d projection_x_coordinate,,,50 -v tasAnom ../../ukcp18-data-factory/fakedata/ukcp18/data/land-prob/uk/25km/rcp85/percentile/tasAnom/mon/latest/tasAnom_rcp85_land-prob_uk_25km_percentile_mon_20001201-20011130.nc ../compliance-check-lib/checklib/test/example_data/tasAnom_rcp85_land-prob_uk_25km_percentile_mon_20001201-20011130.nc" ;
		:NCO = "\"4.5.5\"" ;
data:

 percentile = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 tasAnom = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ; 

 projection_x_coordinate = _ ;

 projection_y_coordinate = _, _ ;
}
